interface d_intf(input logic clk);
  logic d;
  logic rst;
  logic q;
endinterface
